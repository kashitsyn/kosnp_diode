component diode.TcpReceiver

interfaces {
    service : diode.Service
}
