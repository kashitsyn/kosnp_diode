component diode.ConfigurationManager

interfaces {
    dataStorage: diode.DataStorage
}
