component diode.TcpSender

interfaces {
    service : diode.Service
    consumer: diode.Consumer
}
